`ifndef __STATUS_VH__
`define __STATUS_VH__

`define STAT_NORMAL 3'b000
`define STAT_IC_MISS 3'b001
`define STAT_DC_MISS 3'b010
`define STAT_DC_MISS_D 3'b011
`define STAT_DOUBLE_MISS 3'b100
`define STAT_DOUBLE_MISS_D 3'b101

`define COUNT_FINISH 3'd0
`define N_WORDS 3'd4

`endif
