// +FHDR--------------------------------------------------------------------------------------------
// Copyright (c) 2016 Xxx.
// -------------------------------------------------------------------------------------------------
// Filename      : seg_top.v
// Author        : zyy
// Created On    : 2016-05-04 23:41
// Last Modified : 2016-05-04 23:50
// -------------------------------------------------------------------------------------------------
// Svn Info:
//   $Revision::                                                                                $:
//   $Author::                                                                                  $:
//   $Date::                                                                                    $:
//   $HeadURL::                                                                                 $:
// -------------------------------------------------------------------------------------------------
// Description:
//
//
// -FHDR--------------------------------------------------------------------------------------------

module seg_top(
    input clk,
    output [6:0] seg_out,
    output [7:0] seg_ctrl
);

reg [3:0] hex [7:0];

initial begin
    hex[0] <= 4'ha;
    hex[1] <= 4'hb;
    hex[2] <= 4'hc;
    hex[3] <= 4'hd;
    hex[4] <= 4'he;
    hex[5] <= 4'hf;
    hex[6] <= 4'h7;
    hex[7] <= 4'h8;
end

seg_ctrl sc0(
    .clk        (clk        ),
    .hex1       (hex[0]     ),
    .hex2       (hex[1]     ),
    .hex3       (hex[2]     ),
    .hex4       (hex[3]     ),
    .hex5       (hex[4]     ),
    .hex6       (hex[5]     ),
    .hex7       (hex[6]     ),
    .hex8       (hex[7]     ),
    .seg_out    (seg_out    ),
    .seg_ctrl   (seg_ctrl   )
);

endmodule

